--            DO WHAT THE FUCK YOU WANT TO PUBLIC LICENSE
--                    Version 2, December 2004
--
-- Copyright (C) 2004 Sam Hocevar <sam@hocevar.net>
--
-- Everyone is permitted to copy and distribute verbatim or modified
-- copies of this license document, and changing it is allowed as long
-- as the name is changed.
--
--            DO WHAT THE FUCK YOU WANT TO PUBLIC LICENSE
--   TERMS AND CONDITIONS FOR COPYING, DISTRIBUTION AND MODIFICATION
--
--  0. You just DO WHAT THE FUCK YOU WANT TO.
--

-- -- TestBench
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testBenchEvenOdd is
end testBenchEvenOdd;

architecture testEvenOdd of testBenchEvenOdd is

    -- Declare component for TestBench use
    component decideEvenOdd port (
        bit0 : in  std_logic;
        bit1 : in  std_logic;
        bit2 : in  std_logic;
        bit3 : in  std_logic;
        bit4 : in  std_logic;
        bit5 : in  std_logic;
        bit6 : in  std_logic;
        bit7 : in  std_logic;
        bit8 : in  std_logic;
        even:  out std_logic;
        odd:   out std_logic
    ); end component;

    -- Inputs
    signal bit0 : std_logic;
    signal bit1 : std_logic;
    signal bit2 : std_logic;
    signal bit3 : std_logic;
    signal bit4 : std_logic;
    signal bit5 : std_logic;
    signal bit6 : std_logic;
    signal bit7 : std_logic;
    signal bit8 : std_logic;

    -- Outputs
    signal even:  std_logic;
    signal odd:   std_logic;

begin

    -- Creates Even or Odd instance
    deciderInstance: decideEvenOdd port map(
        bit0  => bit0 ,
        bit1  => bit1 ,
        bit2  => bit2 ,
        bit3  => bit3 ,
        bit4  => bit4 ,
        bit5  => bit5 ,
        bit6  => bit6 ,
        bit7  => bit7 ,
        bit8  => bit8 ,
        even  => even,
        odd   => odd
    );

    -- Flips bit 0 every 10 ns
    flippingProcess0: process
        begin loop
            bit0  <= '0';
            wait for 10 ns;
            bit0  <= '1';
            wait for 10 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess0;

    -- Flips bit 1 every 20 ns
    flippingProcess1: process
        begin loop
            bit1  <= '0';
            wait for 20 ns;
            bit1  <= '1';
            wait for 20 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess1;

    -- Flips bit 2 every 40 ns
    flippingProcess2: process
        begin loop
            bit2  <= '0';
            wait for 40 ns;
            bit2  <= '1';
            wait for 40 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess2;

    -- Flips bit 3 every 80 ns
    flippingProcess3: process
        begin loop
            bit3  <= '0';
            wait for 80 ns;
            bit3  <= '1';
            wait for 80 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess3;

    -- Flips bit 4 every 160 ns
    flippingProcess4: process
        begin loop
            bit4  <= '0';
            wait for 160 ns;
            bit4  <= '1';
            wait for 160 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess4;

    -- Flips bit 5 every 320 ns
    flippingProcess5: process
        begin loop
            bit5  <= '0';
            wait for 320 ns;
            bit5  <= '1';
            wait for 320 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess5;

    -- Flips bit 6 every 640 ns
    flippingProcess6: process
        begin loop
            bit6  <= '0';
            wait for 640 ns;
            bit6  <= '1';
            wait for 640 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess6;

    -- Flips bit 7 every 1280 ns
    flippingProcess7: process
        begin loop
            bit7  <= '0';
            wait for 1280 ns;
            bit7  <= '1';
            wait for 1280 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess7;

    -- Flips bit 8 every 2560 ns
    flippingProcess8: process
        begin loop
            bit8  <= '0';
            wait for 2560 ns;
            bit8  <= '1';
            wait for 2560 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess8;
end testEvenOdd;


-- -- Even or Odd decider implementation
library IEEE;
use IEEE.std_logic_1164.all;

entity decideEvenOdd is
    port (
        bit0 : in  std_logic;
        bit1 : in  std_logic;
        bit2 : in  std_logic;
        bit3 : in  std_logic;
        bit4 : in  std_logic;
        bit5 : in  std_logic;
        bit6 : in  std_logic;
        bit7 : in  std_logic;
        bit8 : in  std_logic;
        even:  out std_logic;
        odd:   out std_logic
    );
end decideEvenOdd;

architecture tellMeEvenOdd of decideEvenOdd is
    -- Temporary processing signal (concatenate all bits)
    signal concatenatedBits: std_logic_vector(8 downto 0);
begin
    concatenatedBits <= bit8 & bit7 & bit6 & bit5 & bit4 & bit3 & bit2 & bit1 & bit0;

    -- Truth table for when number is even
    with concatenatedBits select even <=
        '1' when "000000000",
        '0' when "000000001",
        '1' when "000000010",
        '0' when "000000011",
        '1' when "000000100",
        '0' when "000000101",
        '1' when "000000110",
        '0' when "000000111",
        '1' when "000001000",
        '0' when "000001001",
        '1' when "000001010",
        '0' when "000001011",
        '1' when "000001100",
        '0' when "000001101",
        '1' when "000001110",
        '0' when "000001111",
        '1' when "000010000",
        '0' when "000010001",
        '1' when "000010010",
        '0' when "000010011",
        '1' when "000010100",
        '0' when "000010101",
        '1' when "000010110",
        '0' when "000010111",
        '1' when "000011000",
        '0' when "000011001",
        '1' when "000011010",
        '0' when "000011011",
        '1' when "000011100",
        '0' when "000011101",
        '1' when "000011110",
        '0' when "000011111",
        '1' when "000100000",
        '0' when "000100001",
        '1' when "000100010",
        '0' when "000100011",
        '1' when "000100100",
        '0' when "000100101",
        '1' when "000100110",
        '0' when "000100111",
        '1' when "000101000",
        '0' when "000101001",
        '1' when "000101010",
        '0' when "000101011",
        '1' when "000101100",
        '0' when "000101101",
        '1' when "000101110",
        '0' when "000101111",
        '1' when "000110000",
        '0' when "000110001",
        '1' when "000110010",
        '0' when "000110011",
        '1' when "000110100",
        '0' when "000110101",
        '1' when "000110110",
        '0' when "000110111",
        '1' when "000111000",
        '0' when "000111001",
        '1' when "000111010",
        '0' when "000111011",
        '1' when "000111100",
        '0' when "000111101",
        '1' when "000111110",
        '0' when "000111111",
        '1' when "001000000",
        '0' when "001000001",
        '1' when "001000010",
        '0' when "001000011",
        '1' when "001000100",
        '0' when "001000101",
        '1' when "001000110",
        '0' when "001000111",
        '1' when "001001000",
        '0' when "001001001",
        '1' when "001001010",
        '0' when "001001011",
        '1' when "001001100",
        '0' when "001001101",
        '1' when "001001110",
        '0' when "001001111",
        '1' when "001010000",
        '0' when "001010001",
        '1' when "001010010",
        '0' when "001010011",
        '1' when "001010100",
        '0' when "001010101",
        '1' when "001010110",
        '0' when "001010111",
        '1' when "001011000",
        '0' when "001011001",
        '1' when "001011010",
        '0' when "001011011",
        '1' when "001011100",
        '0' when "001011101",
        '1' when "001011110",
        '0' when "001011111",
        '1' when "001100000",
        '0' when "001100001",
        '1' when "001100010",
        '0' when "001100011",
        '1' when "001100100",
        '0' when "001100101",
        '1' when "001100110",
        '0' when "001100111",
        '1' when "001101000",
        '0' when "001101001",
        '1' when "001101010",
        '0' when "001101011",
        '1' when "001101100",
        '0' when "001101101",
        '1' when "001101110",
        '0' when "001101111",
        '1' when "001110000",
        '0' when "001110001",
        '1' when "001110010",
        '0' when "001110011",
        '1' when "001110100",
        '0' when "001110101",
        '1' when "001110110",
        '0' when "001110111",
        '1' when "001111000",
        '0' when "001111001",
        '1' when "001111010",
        '0' when "001111011",
        '1' when "001111100",
        '0' when "001111101",
        '1' when "001111110",
        '0' when "001111111",
        '1' when "010000000",
        '0' when "010000001",
        '1' when "010000010",
        '0' when "010000011",
        '1' when "010000100",
        '0' when "010000101",
        '1' when "010000110",
        '0' when "010000111",
        '1' when "010001000",
        '0' when "010001001",
        '1' when "010001010",
        '0' when "010001011",
        '1' when "010001100",
        '0' when "010001101",
        '1' when "010001110",
        '0' when "010001111",
        '1' when "010010000",
        '0' when "010010001",
        '1' when "010010010",
        '0' when "010010011",
        '1' when "010010100",
        '0' when "010010101",
        '1' when "010010110",
        '0' when "010010111",
        '1' when "010011000",
        '0' when "010011001",
        '1' when "010011010",
        '0' when "010011011",
        '1' when "010011100",
        '0' when "010011101",
        '1' when "010011110",
        '0' when "010011111",
        '1' when "010100000",
        '0' when "010100001",
        '1' when "010100010",
        '0' when "010100011",
        '1' when "010100100",
        '0' when "010100101",
        '1' when "010100110",
        '0' when "010100111",
        '1' when "010101000",
        '0' when "010101001",
        '1' when "010101010",
        '0' when "010101011",
        '1' when "010101100",
        '0' when "010101101",
        '1' when "010101110",
        '0' when "010101111",
        '1' when "010110000",
        '0' when "010110001",
        '1' when "010110010",
        '0' when "010110011",
        '1' when "010110100",
        '0' when "010110101",
        '1' when "010110110",
        '0' when "010110111",
        '1' when "010111000",
        '0' when "010111001",
        '1' when "010111010",
        '0' when "010111011",
        '1' when "010111100",
        '0' when "010111101",
        '1' when "010111110",
        '0' when "010111111",
        '1' when "011000000",
        '0' when "011000001",
        '1' when "011000010",
        '0' when "011000011",
        '1' when "011000100",
        '0' when "011000101",
        '1' when "011000110",
        '0' when "011000111",
        '1' when "011001000",
        '0' when "011001001",
        '1' when "011001010",
        '0' when "011001011",
        '1' when "011001100",
        '0' when "011001101",
        '1' when "011001110",
        '0' when "011001111",
        '1' when "011010000",
        '0' when "011010001",
        '1' when "011010010",
        '0' when "011010011",
        '1' when "011010100",
        '0' when "011010101",
        '1' when "011010110",
        '0' when "011010111",
        '1' when "011011000",
        '0' when "011011001",
        '1' when "011011010",
        '0' when "011011011",
        '1' when "011011100",
        '0' when "011011101",
        '1' when "011011110",
        '0' when "011011111",
        '1' when "011100000",
        '0' when "011100001",
        '1' when "011100010",
        '0' when "011100011",
        '1' when "011100100",
        '0' when "011100101",
        '1' when "011100110",
        '0' when "011100111",
        '1' when "011101000",
        '0' when "011101001",
        '1' when "011101010",
        '0' when "011101011",
        '1' when "011101100",
        '0' when "011101101",
        '1' when "011101110",
        '0' when "011101111",
        '1' when "011110000",
        '0' when "011110001",
        '1' when "011110010",
        '0' when "011110011",
        '1' when "011110100",
        '0' when "011110101",
        '1' when "011110110",
        '0' when "011110111",
        '1' when "011111000",
        '0' when "011111001",
        '1' when "011111010",
        '0' when "011111011",
        '1' when "011111100",
        '0' when "011111101",
        '1' when "011111110",
        '0' when "011111111",
        '1' when "100000000",
        '0' when "100000001",
        '1' when "100000010",
        '0' when "100000011",
        '1' when "100000100",
        '0' when "100000101",
        '1' when "100000110",
        '0' when "100000111",
        '1' when "100001000",
        '0' when "100001001",
        '1' when "100001010",
        '0' when "100001011",
        '1' when "100001100",
        '0' when "100001101",
        '1' when "100001110",
        '0' when "100001111",
        '1' when "100010000",
        '0' when "100010001",
        '1' when "100010010",
        '0' when "100010011",
        '1' when "100010100",
        '0' when "100010101",
        '1' when "100010110",
        '0' when "100010111",
        '1' when "100011000",
        '0' when "100011001",
        '1' when "100011010",
        '0' when "100011011",
        '1' when "100011100",
        '0' when "100011101",
        '1' when "100011110",
        '0' when "100011111",
        '1' when "100100000",
        '0' when "100100001",
        '1' when "100100010",
        '0' when "100100011",
        '1' when "100100100",
        '0' when "100100101",
        '1' when "100100110",
        '0' when "100100111",
        '1' when "100101000",
        '0' when "100101001",
        '1' when "100101010",
        '0' when "100101011",
        '1' when "100101100",
        '0' when "100101101",
        '1' when "100101110",
        '0' when "100101111",
        '1' when "100110000",
        '0' when "100110001",
        '1' when "100110010",
        '0' when "100110011",
        '1' when "100110100",
        '0' when "100110101",
        '1' when "100110110",
        '0' when "100110111",
        '1' when "100111000",
        '0' when "100111001",
        '1' when "100111010",
        '0' when "100111011",
        '1' when "100111100",
        '0' when "100111101",
        '1' when "100111110",
        '0' when "100111111",
        '1' when "101000000",
        '0' when "101000001",
        '1' when "101000010",
        '0' when "101000011",
        '1' when "101000100",
        '0' when "101000101",
        '1' when "101000110",
        '0' when "101000111",
        '1' when "101001000",
        '0' when "101001001",
        '1' when "101001010",
        '0' when "101001011",
        '1' when "101001100",
        '0' when "101001101",
        '1' when "101001110",
        '0' when "101001111",
        '1' when "101010000",
        '0' when "101010001",
        '1' when "101010010",
        '0' when "101010011",
        '1' when "101010100",
        '0' when "101010101",
        '1' when "101010110",
        '0' when "101010111",
        '1' when "101011000",
        '0' when "101011001",
        '1' when "101011010",
        '0' when "101011011",
        '1' when "101011100",
        '0' when "101011101",
        '1' when "101011110",
        '0' when "101011111",
        '1' when "101100000",
        '0' when "101100001",
        '1' when "101100010",
        '0' when "101100011",
        '1' when "101100100",
        '0' when "101100101",
        '1' when "101100110",
        '0' when "101100111",
        '1' when "101101000",
        '0' when "101101001",
        '1' when "101101010",
        '0' when "101101011",
        '1' when "101101100",
        '0' when "101101101",
        '1' when "101101110",
        '0' when "101101111",
        '1' when "101110000",
        '0' when "101110001",
        '1' when "101110010",
        '0' when "101110011",
        '1' when "101110100",
        '0' when "101110101",
        '1' when "101110110",
        '0' when "101110111",
        '1' when "101111000",
        '0' when "101111001",
        '1' when "101111010",
        '0' when "101111011",
        '1' when "101111100",
        '0' when "101111101",
        '1' when "101111110",
        '0' when "101111111",
        '1' when "110000000",
        '0' when "110000001",
        '1' when "110000010",
        '0' when "110000011",
        '1' when "110000100",
        '0' when "110000101",
        '1' when "110000110",
        '0' when "110000111",
        '1' when "110001000",
        '0' when "110001001",
        '1' when "110001010",
        '0' when "110001011",
        '1' when "110001100",
        '0' when "110001101",
        '1' when "110001110",
        '0' when "110001111",
        '1' when "110010000",
        '0' when "110010001",
        '1' when "110010010",
        '0' when "110010011",
        '1' when "110010100",
        '0' when "110010101",
        '1' when "110010110",
        '0' when "110010111",
        '1' when "110011000",
        '0' when "110011001",
        '1' when "110011010",
        '0' when "110011011",
        '1' when "110011100",
        '0' when "110011101",
        '1' when "110011110",
        '0' when "110011111",
        '1' when "110100000",
        '0' when "110100001",
        '1' when "110100010",
        '0' when "110100011",
        '1' when "110100100",
        '0' when "110100101",
        '1' when "110100110",
        '0' when "110100111",
        '1' when "110101000",
        '0' when "110101001",
        '1' when "110101010",
        '0' when "110101011",
        '1' when "110101100",
        '0' when "110101101",
        '1' when "110101110",
        '0' when "110101111",
        '1' when "110110000",
        '0' when "110110001",
        '1' when "110110010",
        '0' when "110110011",
        '1' when "110110100",
        '0' when "110110101",
        '1' when "110110110",
        '0' when "110110111",
        '1' when "110111000",
        '0' when "110111001",
        '1' when "110111010",
        '0' when "110111011",
        '1' when "110111100",
        '0' when "110111101",
        '1' when "110111110",
        '0' when "110111111",
        '1' when "111000000",
        '0' when "111000001",
        '1' when "111000010",
        '0' when "111000011",
        '1' when "111000100",
        '0' when "111000101",
        '1' when "111000110",
        '0' when "111000111",
        '1' when "111001000",
        '0' when "111001001",
        '1' when "111001010",
        '0' when "111001011",
        '1' when "111001100",
        '0' when "111001101",
        '1' when "111001110",
        '0' when "111001111",
        '1' when "111010000",
        '0' when "111010001",
        '1' when "111010010",
        '0' when "111010011",
        '1' when "111010100",
        '0' when "111010101",
        '1' when "111010110",
        '0' when "111010111",
        '1' when "111011000",
        '0' when "111011001",
        '1' when "111011010",
        '0' when "111011011",
        '1' when "111011100",
        '0' when "111011101",
        '1' when "111011110",
        '0' when "111011111",
        '1' when "111100000",
        '0' when "111100001",
        '1' when "111100010",
        '0' when "111100011",
        '1' when "111100100",
        '0' when "111100101",
        '1' when "111100110",
        '0' when "111100111",
        '1' when "111101000",
        '0' when "111101001",
        '1' when "111101010",
        '0' when "111101011",
        '1' when "111101100",
        '0' when "111101101",
        '1' when "111101110",
        '0' when "111101111",
        '1' when "111110000",
        '0' when "111110001",
        '1' when "111110010",
        '0' when "111110011",
        '1' when "111110100",
        '0' when "111110101",
        '1' when "111110110",
        '0' when "111110111",
        '1' when "111111000",
        '0' when "111111001",
        '1' when "111111010",
        '0' when "111111011",
        '1' when "111111100",
        '0' when "111111101",
        '1' when "111111110",
        '0' when "111111111",
        '0' when others;

    -- Truth table for when number is odd
    with concatenatedBits select odd <=
        '0' when "000000000",
        '1' when "000000001",
        '0' when "000000010",
        '1' when "000000011",
        '0' when "000000100",
        '1' when "000000101",
        '0' when "000000110",
        '1' when "000000111",
        '0' when "000001000",
        '1' when "000001001",
        '0' when "000001010",
        '1' when "000001011",
        '0' when "000001100",
        '1' when "000001101",
        '0' when "000001110",
        '1' when "000001111",
        '0' when "000010000",
        '1' when "000010001",
        '0' when "000010010",
        '1' when "000010011",
        '0' when "000010100",
        '1' when "000010101",
        '0' when "000010110",
        '1' when "000010111",
        '0' when "000011000",
        '1' when "000011001",
        '0' when "000011010",
        '1' when "000011011",
        '0' when "000011100",
        '1' when "000011101",
        '0' when "000011110",
        '1' when "000011111",
        '0' when "000100000",
        '1' when "000100001",
        '0' when "000100010",
        '1' when "000100011",
        '0' when "000100100",
        '1' when "000100101",
        '0' when "000100110",
        '1' when "000100111",
        '0' when "000101000",
        '1' when "000101001",
        '0' when "000101010",
        '1' when "000101011",
        '0' when "000101100",
        '1' when "000101101",
        '0' when "000101110",
        '1' when "000101111",
        '0' when "000110000",
        '1' when "000110001",
        '0' when "000110010",
        '1' when "000110011",
        '0' when "000110100",
        '1' when "000110101",
        '0' when "000110110",
        '1' when "000110111",
        '0' when "000111000",
        '1' when "000111001",
        '0' when "000111010",
        '1' when "000111011",
        '0' when "000111100",
        '1' when "000111101",
        '0' when "000111110",
        '1' when "000111111",
        '0' when "001000000",
        '1' when "001000001",
        '0' when "001000010",
        '1' when "001000011",
        '0' when "001000100",
        '1' when "001000101",
        '0' when "001000110",
        '1' when "001000111",
        '0' when "001001000",
        '1' when "001001001",
        '0' when "001001010",
        '1' when "001001011",
        '0' when "001001100",
        '1' when "001001101",
        '0' when "001001110",
        '1' when "001001111",
        '0' when "001010000",
        '1' when "001010001",
        '0' when "001010010",
        '1' when "001010011",
        '0' when "001010100",
        '1' when "001010101",
        '0' when "001010110",
        '1' when "001010111",
        '0' when "001011000",
        '1' when "001011001",
        '0' when "001011010",
        '1' when "001011011",
        '0' when "001011100",
        '1' when "001011101",
        '0' when "001011110",
        '1' when "001011111",
        '0' when "001100000",
        '1' when "001100001",
        '0' when "001100010",
        '1' when "001100011",
        '0' when "001100100",
        '1' when "001100101",
        '0' when "001100110",
        '1' when "001100111",
        '0' when "001101000",
        '1' when "001101001",
        '0' when "001101010",
        '1' when "001101011",
        '0' when "001101100",
        '1' when "001101101",
        '0' when "001101110",
        '1' when "001101111",
        '0' when "001110000",
        '1' when "001110001",
        '0' when "001110010",
        '1' when "001110011",
        '0' when "001110100",
        '1' when "001110101",
        '0' when "001110110",
        '1' when "001110111",
        '0' when "001111000",
        '1' when "001111001",
        '0' when "001111010",
        '1' when "001111011",
        '0' when "001111100",
        '1' when "001111101",
        '0' when "001111110",
        '1' when "001111111",
        '0' when "010000000",
        '1' when "010000001",
        '0' when "010000010",
        '1' when "010000011",
        '0' when "010000100",
        '1' when "010000101",
        '0' when "010000110",
        '1' when "010000111",
        '0' when "010001000",
        '1' when "010001001",
        '0' when "010001010",
        '1' when "010001011",
        '0' when "010001100",
        '1' when "010001101",
        '0' when "010001110",
        '1' when "010001111",
        '0' when "010010000",
        '1' when "010010001",
        '0' when "010010010",
        '1' when "010010011",
        '0' when "010010100",
        '1' when "010010101",
        '0' when "010010110",
        '1' when "010010111",
        '0' when "010011000",
        '1' when "010011001",
        '0' when "010011010",
        '1' when "010011011",
        '0' when "010011100",
        '1' when "010011101",
        '0' when "010011110",
        '1' when "010011111",
        '0' when "010100000",
        '1' when "010100001",
        '0' when "010100010",
        '1' when "010100011",
        '0' when "010100100",
        '1' when "010100101",
        '0' when "010100110",
        '1' when "010100111",
        '0' when "010101000",
        '1' when "010101001",
        '0' when "010101010",
        '1' when "010101011",
        '0' when "010101100",
        '1' when "010101101",
        '0' when "010101110",
        '1' when "010101111",
        '0' when "010110000",
        '1' when "010110001",
        '0' when "010110010",
        '1' when "010110011",
        '0' when "010110100",
        '1' when "010110101",
        '0' when "010110110",
        '1' when "010110111",
        '0' when "010111000",
        '1' when "010111001",
        '0' when "010111010",
        '1' when "010111011",
        '0' when "010111100",
        '1' when "010111101",
        '0' when "010111110",
        '1' when "010111111",
        '0' when "011000000",
        '1' when "011000001",
        '0' when "011000010",
        '1' when "011000011",
        '0' when "011000100",
        '1' when "011000101",
        '0' when "011000110",
        '1' when "011000111",
        '0' when "011001000",
        '1' when "011001001",
        '0' when "011001010",
        '1' when "011001011",
        '0' when "011001100",
        '1' when "011001101",
        '0' when "011001110",
        '1' when "011001111",
        '0' when "011010000",
        '1' when "011010001",
        '0' when "011010010",
        '1' when "011010011",
        '0' when "011010100",
        '1' when "011010101",
        '0' when "011010110",
        '1' when "011010111",
        '0' when "011011000",
        '1' when "011011001",
        '0' when "011011010",
        '1' when "011011011",
        '0' when "011011100",
        '1' when "011011101",
        '0' when "011011110",
        '1' when "011011111",
        '0' when "011100000",
        '1' when "011100001",
        '0' when "011100010",
        '1' when "011100011",
        '0' when "011100100",
        '1' when "011100101",
        '0' when "011100110",
        '1' when "011100111",
        '0' when "011101000",
        '1' when "011101001",
        '0' when "011101010",
        '1' when "011101011",
        '0' when "011101100",
        '1' when "011101101",
        '0' when "011101110",
        '1' when "011101111",
        '0' when "011110000",
        '1' when "011110001",
        '0' when "011110010",
        '1' when "011110011",
        '0' when "011110100",
        '1' when "011110101",
        '0' when "011110110",
        '1' when "011110111",
        '0' when "011111000",
        '1' when "011111001",
        '0' when "011111010",
        '1' when "011111011",
        '0' when "011111100",
        '1' when "011111101",
        '0' when "011111110",
        '1' when "011111111",
        '0' when "100000000",
        '1' when "100000001",
        '0' when "100000010",
        '1' when "100000011",
        '0' when "100000100",
        '1' when "100000101",
        '0' when "100000110",
        '1' when "100000111",
        '0' when "100001000",
        '1' when "100001001",
        '0' when "100001010",
        '1' when "100001011",
        '0' when "100001100",
        '1' when "100001101",
        '0' when "100001110",
        '1' when "100001111",
        '0' when "100010000",
        '1' when "100010001",
        '0' when "100010010",
        '1' when "100010011",
        '0' when "100010100",
        '1' when "100010101",
        '0' when "100010110",
        '1' when "100010111",
        '0' when "100011000",
        '1' when "100011001",
        '0' when "100011010",
        '1' when "100011011",
        '0' when "100011100",
        '1' when "100011101",
        '0' when "100011110",
        '1' when "100011111",
        '0' when "100100000",
        '1' when "100100001",
        '0' when "100100010",
        '1' when "100100011",
        '0' when "100100100",
        '1' when "100100101",
        '0' when "100100110",
        '1' when "100100111",
        '0' when "100101000",
        '1' when "100101001",
        '0' when "100101010",
        '1' when "100101011",
        '0' when "100101100",
        '1' when "100101101",
        '0' when "100101110",
        '1' when "100101111",
        '0' when "100110000",
        '1' when "100110001",
        '0' when "100110010",
        '1' when "100110011",
        '0' when "100110100",
        '1' when "100110101",
        '0' when "100110110",
        '1' when "100110111",
        '0' when "100111000",
        '1' when "100111001",
        '0' when "100111010",
        '1' when "100111011",
        '0' when "100111100",
        '1' when "100111101",
        '0' when "100111110",
        '1' when "100111111",
        '0' when "101000000",
        '1' when "101000001",
        '0' when "101000010",
        '1' when "101000011",
        '0' when "101000100",
        '1' when "101000101",
        '0' when "101000110",
        '1' when "101000111",
        '0' when "101001000",
        '1' when "101001001",
        '0' when "101001010",
        '1' when "101001011",
        '0' when "101001100",
        '1' when "101001101",
        '0' when "101001110",
        '1' when "101001111",
        '0' when "101010000",
        '1' when "101010001",
        '0' when "101010010",
        '1' when "101010011",
        '0' when "101010100",
        '1' when "101010101",
        '0' when "101010110",
        '1' when "101010111",
        '0' when "101011000",
        '1' when "101011001",
        '0' when "101011010",
        '1' when "101011011",
        '0' when "101011100",
        '1' when "101011101",
        '0' when "101011110",
        '1' when "101011111",
        '0' when "101100000",
        '1' when "101100001",
        '0' when "101100010",
        '1' when "101100011",
        '0' when "101100100",
        '1' when "101100101",
        '0' when "101100110",
        '1' when "101100111",
        '0' when "101101000",
        '1' when "101101001",
        '0' when "101101010",
        '1' when "101101011",
        '0' when "101101100",
        '1' when "101101101",
        '0' when "101101110",
        '1' when "101101111",
        '0' when "101110000",
        '1' when "101110001",
        '0' when "101110010",
        '1' when "101110011",
        '0' when "101110100",
        '1' when "101110101",
        '0' when "101110110",
        '1' when "101110111",
        '0' when "101111000",
        '1' when "101111001",
        '0' when "101111010",
        '1' when "101111011",
        '0' when "101111100",
        '1' when "101111101",
        '0' when "101111110",
        '1' when "101111111",
        '0' when "110000000",
        '1' when "110000001",
        '0' when "110000010",
        '1' when "110000011",
        '0' when "110000100",
        '1' when "110000101",
        '0' when "110000110",
        '1' when "110000111",
        '0' when "110001000",
        '1' when "110001001",
        '0' when "110001010",
        '1' when "110001011",
        '0' when "110001100",
        '1' when "110001101",
        '0' when "110001110",
        '1' when "110001111",
        '0' when "110010000",
        '1' when "110010001",
        '0' when "110010010",
        '1' when "110010011",
        '0' when "110010100",
        '1' when "110010101",
        '0' when "110010110",
        '1' when "110010111",
        '0' when "110011000",
        '1' when "110011001",
        '0' when "110011010",
        '1' when "110011011",
        '0' when "110011100",
        '1' when "110011101",
        '0' when "110011110",
        '1' when "110011111",
        '0' when "110100000",
        '1' when "110100001",
        '0' when "110100010",
        '1' when "110100011",
        '0' when "110100100",
        '1' when "110100101",
        '0' when "110100110",
        '1' when "110100111",
        '0' when "110101000",
        '1' when "110101001",
        '0' when "110101010",
        '1' when "110101011",
        '0' when "110101100",
        '1' when "110101101",
        '0' when "110101110",
        '1' when "110101111",
        '0' when "110110000",
        '1' when "110110001",
        '0' when "110110010",
        '1' when "110110011",
        '0' when "110110100",
        '1' when "110110101",
        '0' when "110110110",
        '1' when "110110111",
        '0' when "110111000",
        '1' when "110111001",
        '0' when "110111010",
        '1' when "110111011",
        '0' when "110111100",
        '1' when "110111101",
        '0' when "110111110",
        '1' when "110111111",
        '0' when "111000000",
        '1' when "111000001",
        '0' when "111000010",
        '1' when "111000011",
        '0' when "111000100",
        '1' when "111000101",
        '0' when "111000110",
        '1' when "111000111",
        '0' when "111001000",
        '1' when "111001001",
        '0' when "111001010",
        '1' when "111001011",
        '0' when "111001100",
        '1' when "111001101",
        '0' when "111001110",
        '1' when "111001111",
        '0' when "111010000",
        '1' when "111010001",
        '0' when "111010010",
        '1' when "111010011",
        '0' when "111010100",
        '1' when "111010101",
        '0' when "111010110",
        '1' when "111010111",
        '0' when "111011000",
        '1' when "111011001",
        '0' when "111011010",
        '1' when "111011011",
        '0' when "111011100",
        '1' when "111011101",
        '0' when "111011110",
        '1' when "111011111",
        '0' when "111100000",
        '1' when "111100001",
        '0' when "111100010",
        '1' when "111100011",
        '0' when "111100100",
        '1' when "111100101",
        '0' when "111100110",
        '1' when "111100111",
        '0' when "111101000",
        '1' when "111101001",
        '0' when "111101010",
        '1' when "111101011",
        '0' when "111101100",
        '1' when "111101101",
        '0' when "111101110",
        '1' when "111101111",
        '0' when "111110000",
        '1' when "111110001",
        '0' when "111110010",
        '1' when "111110011",
        '0' when "111110100",
        '1' when "111110101",
        '0' when "111110110",
        '1' when "111110111",
        '0' when "111111000",
        '1' when "111111001",
        '0' when "111111010",
        '1' when "111111011",
        '0' when "111111100",
        '1' when "111111101",
        '0' when "111111110",
        '1' when "111111111",
        '0' when others;
end tellMeEvenOdd;

-- Thanks for using my library, hope you have memory for it!!
-- (The speeds are theoretically massive, memory is not an issue)