--            DO WHAT THE FUCK YOU WANT TO PUBLIC LICENSE
--                    Version 2, December 2004
--
-- Copyright (C) 2004 Sam Hocevar <sam@hocevar.net>
--
-- Everyone is permitted to copy and distribute verbatim or modified
-- copies of this license document, and changing it is allowed as long
-- as the name is changed.
--
--            DO WHAT THE FUCK YOU WANT TO PUBLIC LICENSE
--   TERMS AND CONDITIONS FOR COPYING, DISTRIBUTION AND MODIFICATION
--
--  0. You just DO WHAT THE FUCK YOU WANT TO.
--

-- -- TestBench
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testBenchEvenOdd is
end testBenchEvenOdd;

architecture testEvenOdd of testBenchEvenOdd is

    -- Declare component for TestBench use
    component decideEvenOdd port (
        bit0 : in  std_logic;
        bit1 : in  std_logic;
        bit2 : in  std_logic;
        bit3 : in  std_logic;
        bit4 : in  std_logic;
        bit5 : in  std_logic;
        bit6 : in  std_logic;
        bit7 : in  std_logic;
        bit8 : in  std_logic;
        bit9 : in  std_logic;
        even:  out std_logic;
        odd:   out std_logic
    ); end component;

    -- Inputs
    signal bit0 : std_logic;
    signal bit1 : std_logic;
    signal bit2 : std_logic;
    signal bit3 : std_logic;
    signal bit4 : std_logic;
    signal bit5 : std_logic;
    signal bit6 : std_logic;
    signal bit7 : std_logic;
    signal bit8 : std_logic;
    signal bit9 : std_logic;

    -- Outputs
    signal even:  std_logic;
    signal odd:   std_logic;

begin

    -- Creates Even or Odd instance
    deciderInstance: decideEvenOdd port map(
        bit0  => bit0 ,
        bit1  => bit1 ,
        bit2  => bit2 ,
        bit3  => bit3 ,
        bit4  => bit4 ,
        bit5  => bit5 ,
        bit6  => bit6 ,
        bit7  => bit7 ,
        bit8  => bit8 ,
        bit9  => bit9 ,
        even  => even,
        odd   => odd
    );

    -- Flips bit 0 every 10 ns
    flippingProcess0: process
        begin loop
            bit0  <= '0';
            wait for 10 ns;
            bit0  <= '1';
            wait for 10 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess0;

    -- Flips bit 1 every 20 ns
    flippingProcess1: process
        begin loop
            bit1  <= '0';
            wait for 20 ns;
            bit1  <= '1';
            wait for 20 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess1;

    -- Flips bit 2 every 40 ns
    flippingProcess2: process
        begin loop
            bit2  <= '0';
            wait for 40 ns;
            bit2  <= '1';
            wait for 40 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess2;

    -- Flips bit 3 every 80 ns
    flippingProcess3: process
        begin loop
            bit3  <= '0';
            wait for 80 ns;
            bit3  <= '1';
            wait for 80 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess3;

    -- Flips bit 4 every 160 ns
    flippingProcess4: process
        begin loop
            bit4  <= '0';
            wait for 160 ns;
            bit4  <= '1';
            wait for 160 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess4;

    -- Flips bit 5 every 320 ns
    flippingProcess5: process
        begin loop
            bit5  <= '0';
            wait for 320 ns;
            bit5  <= '1';
            wait for 320 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess5;

    -- Flips bit 6 every 640 ns
    flippingProcess6: process
        begin loop
            bit6  <= '0';
            wait for 640 ns;
            bit6  <= '1';
            wait for 640 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess6;

    -- Flips bit 7 every 1280 ns
    flippingProcess7: process
        begin loop
            bit7  <= '0';
            wait for 1280 ns;
            bit7  <= '1';
            wait for 1280 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess7;

    -- Flips bit 8 every 2560 ns
    flippingProcess8: process
        begin loop
            bit8  <= '0';
            wait for 2560 ns;
            bit8  <= '1';
            wait for 2560 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess8;

    -- Flips bit 9 every 5120 ns
    flippingProcess9: process
        begin loop
            bit9  <= '0';
            wait for 5120 ns;
            bit9  <= '1';
            wait for 5120 ns;
            if NOW > 3200 ns then wait; end if;
        end loop;
    end process flippingProcess9;
end testEvenOdd;


-- -- Even or Odd decider implementation
library IEEE;
use IEEE.std_logic_1164.all;

entity decideEvenOdd is
    port (
        bit0 : in  std_logic;
        bit1 : in  std_logic;
        bit2 : in  std_logic;
        bit3 : in  std_logic;
        bit4 : in  std_logic;
        bit5 : in  std_logic;
        bit6 : in  std_logic;
        bit7 : in  std_logic;
        bit8 : in  std_logic;
        bit9 : in  std_logic;
        even:  out std_logic;
        odd:   out std_logic
    );
end decideEvenOdd;

architecture tellMeEvenOdd of decideEvenOdd is
    -- Temporary processing signal (concatenate all bits)
    signal concatenatedBits: std_logic_vector(9 downto 0);
begin
    concatenatedBits <= bit9 & bit8 & bit7 & bit6 & bit5 & bit4 & bit3 & bit2 & bit1 & bit0;

    -- Truth table for when number is even
    with concatenatedBits select even <=
        '1' when "0000000000",
        '0' when "0000000001",
        '1' when "0000000010",
        '0' when "0000000011",
        '1' when "0000000100",
        '0' when "0000000101",
        '1' when "0000000110",
        '0' when "0000000111",
        '1' when "0000001000",
        '0' when "0000001001",
        '1' when "0000001010",
        '0' when "0000001011",
        '1' when "0000001100",
        '0' when "0000001101",
        '1' when "0000001110",
        '0' when "0000001111",
        '1' when "0000010000",
        '0' when "0000010001",
        '1' when "0000010010",
        '0' when "0000010011",
        '1' when "0000010100",
        '0' when "0000010101",
        '1' when "0000010110",
        '0' when "0000010111",
        '1' when "0000011000",
        '0' when "0000011001",
        '1' when "0000011010",
        '0' when "0000011011",
        '1' when "0000011100",
        '0' when "0000011101",
        '1' when "0000011110",
        '0' when "0000011111",
        '1' when "0000100000",
        '0' when "0000100001",
        '1' when "0000100010",
        '0' when "0000100011",
        '1' when "0000100100",
        '0' when "0000100101",
        '1' when "0000100110",
        '0' when "0000100111",
        '1' when "0000101000",
        '0' when "0000101001",
        '1' when "0000101010",
        '0' when "0000101011",
        '1' when "0000101100",
        '0' when "0000101101",
        '1' when "0000101110",
        '0' when "0000101111",
        '1' when "0000110000",
        '0' when "0000110001",
        '1' when "0000110010",
        '0' when "0000110011",
        '1' when "0000110100",
        '0' when "0000110101",
        '1' when "0000110110",
        '0' when "0000110111",
        '1' when "0000111000",
        '0' when "0000111001",
        '1' when "0000111010",
        '0' when "0000111011",
        '1' when "0000111100",
        '0' when "0000111101",
        '1' when "0000111110",
        '0' when "0000111111",
        '1' when "0001000000",
        '0' when "0001000001",
        '1' when "0001000010",
        '0' when "0001000011",
        '1' when "0001000100",
        '0' when "0001000101",
        '1' when "0001000110",
        '0' when "0001000111",
        '1' when "0001001000",
        '0' when "0001001001",
        '1' when "0001001010",
        '0' when "0001001011",
        '1' when "0001001100",
        '0' when "0001001101",
        '1' when "0001001110",
        '0' when "0001001111",
        '1' when "0001010000",
        '0' when "0001010001",
        '1' when "0001010010",
        '0' when "0001010011",
        '1' when "0001010100",
        '0' when "0001010101",
        '1' when "0001010110",
        '0' when "0001010111",
        '1' when "0001011000",
        '0' when "0001011001",
        '1' when "0001011010",
        '0' when "0001011011",
        '1' when "0001011100",
        '0' when "0001011101",
        '1' when "0001011110",
        '0' when "0001011111",
        '1' when "0001100000",
        '0' when "0001100001",
        '1' when "0001100010",
        '0' when "0001100011",
        '1' when "0001100100",
        '0' when "0001100101",
        '1' when "0001100110",
        '0' when "0001100111",
        '1' when "0001101000",
        '0' when "0001101001",
        '1' when "0001101010",
        '0' when "0001101011",
        '1' when "0001101100",
        '0' when "0001101101",
        '1' when "0001101110",
        '0' when "0001101111",
        '1' when "0001110000",
        '0' when "0001110001",
        '1' when "0001110010",
        '0' when "0001110011",
        '1' when "0001110100",
        '0' when "0001110101",
        '1' when "0001110110",
        '0' when "0001110111",
        '1' when "0001111000",
        '0' when "0001111001",
        '1' when "0001111010",
        '0' when "0001111011",
        '1' when "0001111100",
        '0' when "0001111101",
        '1' when "0001111110",
        '0' when "0001111111",
        '1' when "0010000000",
        '0' when "0010000001",
        '1' when "0010000010",
        '0' when "0010000011",
        '1' when "0010000100",
        '0' when "0010000101",
        '1' when "0010000110",
        '0' when "0010000111",
        '1' when "0010001000",
        '0' when "0010001001",
        '1' when "0010001010",
        '0' when "0010001011",
        '1' when "0010001100",
        '0' when "0010001101",
        '1' when "0010001110",
        '0' when "0010001111",
        '1' when "0010010000",
        '0' when "0010010001",
        '1' when "0010010010",
        '0' when "0010010011",
        '1' when "0010010100",
        '0' when "0010010101",
        '1' when "0010010110",
        '0' when "0010010111",
        '1' when "0010011000",
        '0' when "0010011001",
        '1' when "0010011010",
        '0' when "0010011011",
        '1' when "0010011100",
        '0' when "0010011101",
        '1' when "0010011110",
        '0' when "0010011111",
        '1' when "0010100000",
        '0' when "0010100001",
        '1' when "0010100010",
        '0' when "0010100011",
        '1' when "0010100100",
        '0' when "0010100101",
        '1' when "0010100110",
        '0' when "0010100111",
        '1' when "0010101000",
        '0' when "0010101001",
        '1' when "0010101010",
        '0' when "0010101011",
        '1' when "0010101100",
        '0' when "0010101101",
        '1' when "0010101110",
        '0' when "0010101111",
        '1' when "0010110000",
        '0' when "0010110001",
        '1' when "0010110010",
        '0' when "0010110011",
        '1' when "0010110100",
        '0' when "0010110101",
        '1' when "0010110110",
        '0' when "0010110111",
        '1' when "0010111000",
        '0' when "0010111001",
        '1' when "0010111010",
        '0' when "0010111011",
        '1' when "0010111100",
        '0' when "0010111101",
        '1' when "0010111110",
        '0' when "0010111111",
        '1' when "0011000000",
        '0' when "0011000001",
        '1' when "0011000010",
        '0' when "0011000011",
        '1' when "0011000100",
        '0' when "0011000101",
        '1' when "0011000110",
        '0' when "0011000111",
        '1' when "0011001000",
        '0' when "0011001001",
        '1' when "0011001010",
        '0' when "0011001011",
        '1' when "0011001100",
        '0' when "0011001101",
        '1' when "0011001110",
        '0' when "0011001111",
        '1' when "0011010000",
        '0' when "0011010001",
        '1' when "0011010010",
        '0' when "0011010011",
        '1' when "0011010100",
        '0' when "0011010101",
        '1' when "0011010110",
        '0' when "0011010111",
        '1' when "0011011000",
        '0' when "0011011001",
        '1' when "0011011010",
        '0' when "0011011011",
        '1' when "0011011100",
        '0' when "0011011101",
        '1' when "0011011110",
        '0' when "0011011111",
        '1' when "0011100000",
        '0' when "0011100001",
        '1' when "0011100010",
        '0' when "0011100011",
        '1' when "0011100100",
        '0' when "0011100101",
        '1' when "0011100110",
        '0' when "0011100111",
        '1' when "0011101000",
        '0' when "0011101001",
        '1' when "0011101010",
        '0' when "0011101011",
        '1' when "0011101100",
        '0' when "0011101101",
        '1' when "0011101110",
        '0' when "0011101111",
        '1' when "0011110000",
        '0' when "0011110001",
        '1' when "0011110010",
        '0' when "0011110011",
        '1' when "0011110100",
        '0' when "0011110101",
        '1' when "0011110110",
        '0' when "0011110111",
        '1' when "0011111000",
        '0' when "0011111001",
        '1' when "0011111010",
        '0' when "0011111011",
        '1' when "0011111100",
        '0' when "0011111101",
        '1' when "0011111110",
        '0' when "0011111111",
        '1' when "0100000000",
        '0' when "0100000001",
        '1' when "0100000010",
        '0' when "0100000011",
        '1' when "0100000100",
        '0' when "0100000101",
        '1' when "0100000110",
        '0' when "0100000111",
        '1' when "0100001000",
        '0' when "0100001001",
        '1' when "0100001010",
        '0' when "0100001011",
        '1' when "0100001100",
        '0' when "0100001101",
        '1' when "0100001110",
        '0' when "0100001111",
        '1' when "0100010000",
        '0' when "0100010001",
        '1' when "0100010010",
        '0' when "0100010011",
        '1' when "0100010100",
        '0' when "0100010101",
        '1' when "0100010110",
        '0' when "0100010111",
        '1' when "0100011000",
        '0' when "0100011001",
        '1' when "0100011010",
        '0' when "0100011011",
        '1' when "0100011100",
        '0' when "0100011101",
        '1' when "0100011110",
        '0' when "0100011111",
        '1' when "0100100000",
        '0' when "0100100001",
        '1' when "0100100010",
        '0' when "0100100011",
        '1' when "0100100100",
        '0' when "0100100101",
        '1' when "0100100110",
        '0' when "0100100111",
        '1' when "0100101000",
        '0' when "0100101001",
        '1' when "0100101010",
        '0' when "0100101011",
        '1' when "0100101100",
        '0' when "0100101101",
        '1' when "0100101110",
        '0' when "0100101111",
        '1' when "0100110000",
        '0' when "0100110001",
        '1' when "0100110010",
        '0' when "0100110011",
        '1' when "0100110100",
        '0' when "0100110101",
        '1' when "0100110110",
        '0' when "0100110111",
        '1' when "0100111000",
        '0' when "0100111001",
        '1' when "0100111010",
        '0' when "0100111011",
        '1' when "0100111100",
        '0' when "0100111101",
        '1' when "0100111110",
        '0' when "0100111111",
        '1' when "0101000000",
        '0' when "0101000001",
        '1' when "0101000010",
        '0' when "0101000011",
        '1' when "0101000100",
        '0' when "0101000101",
        '1' when "0101000110",
        '0' when "0101000111",
        '1' when "0101001000",
        '0' when "0101001001",
        '1' when "0101001010",
        '0' when "0101001011",
        '1' when "0101001100",
        '0' when "0101001101",
        '1' when "0101001110",
        '0' when "0101001111",
        '1' when "0101010000",
        '0' when "0101010001",
        '1' when "0101010010",
        '0' when "0101010011",
        '1' when "0101010100",
        '0' when "0101010101",
        '1' when "0101010110",
        '0' when "0101010111",
        '1' when "0101011000",
        '0' when "0101011001",
        '1' when "0101011010",
        '0' when "0101011011",
        '1' when "0101011100",
        '0' when "0101011101",
        '1' when "0101011110",
        '0' when "0101011111",
        '1' when "0101100000",
        '0' when "0101100001",
        '1' when "0101100010",
        '0' when "0101100011",
        '1' when "0101100100",
        '0' when "0101100101",
        '1' when "0101100110",
        '0' when "0101100111",
        '1' when "0101101000",
        '0' when "0101101001",
        '1' when "0101101010",
        '0' when "0101101011",
        '1' when "0101101100",
        '0' when "0101101101",
        '1' when "0101101110",
        '0' when "0101101111",
        '1' when "0101110000",
        '0' when "0101110001",
        '1' when "0101110010",
        '0' when "0101110011",
        '1' when "0101110100",
        '0' when "0101110101",
        '1' when "0101110110",
        '0' when "0101110111",
        '1' when "0101111000",
        '0' when "0101111001",
        '1' when "0101111010",
        '0' when "0101111011",
        '1' when "0101111100",
        '0' when "0101111101",
        '1' when "0101111110",
        '0' when "0101111111",
        '1' when "0110000000",
        '0' when "0110000001",
        '1' when "0110000010",
        '0' when "0110000011",
        '1' when "0110000100",
        '0' when "0110000101",
        '1' when "0110000110",
        '0' when "0110000111",
        '1' when "0110001000",
        '0' when "0110001001",
        '1' when "0110001010",
        '0' when "0110001011",
        '1' when "0110001100",
        '0' when "0110001101",
        '1' when "0110001110",
        '0' when "0110001111",
        '1' when "0110010000",
        '0' when "0110010001",
        '1' when "0110010010",
        '0' when "0110010011",
        '1' when "0110010100",
        '0' when "0110010101",
        '1' when "0110010110",
        '0' when "0110010111",
        '1' when "0110011000",
        '0' when "0110011001",
        '1' when "0110011010",
        '0' when "0110011011",
        '1' when "0110011100",
        '0' when "0110011101",
        '1' when "0110011110",
        '0' when "0110011111",
        '1' when "0110100000",
        '0' when "0110100001",
        '1' when "0110100010",
        '0' when "0110100011",
        '1' when "0110100100",
        '0' when "0110100101",
        '1' when "0110100110",
        '0' when "0110100111",
        '1' when "0110101000",
        '0' when "0110101001",
        '1' when "0110101010",
        '0' when "0110101011",
        '1' when "0110101100",
        '0' when "0110101101",
        '1' when "0110101110",
        '0' when "0110101111",
        '1' when "0110110000",
        '0' when "0110110001",
        '1' when "0110110010",
        '0' when "0110110011",
        '1' when "0110110100",
        '0' when "0110110101",
        '1' when "0110110110",
        '0' when "0110110111",
        '1' when "0110111000",
        '0' when "0110111001",
        '1' when "0110111010",
        '0' when "0110111011",
        '1' when "0110111100",
        '0' when "0110111101",
        '1' when "0110111110",
        '0' when "0110111111",
        '1' when "0111000000",
        '0' when "0111000001",
        '1' when "0111000010",
        '0' when "0111000011",
        '1' when "0111000100",
        '0' when "0111000101",
        '1' when "0111000110",
        '0' when "0111000111",
        '1' when "0111001000",
        '0' when "0111001001",
        '1' when "0111001010",
        '0' when "0111001011",
        '1' when "0111001100",
        '0' when "0111001101",
        '1' when "0111001110",
        '0' when "0111001111",
        '1' when "0111010000",
        '0' when "0111010001",
        '1' when "0111010010",
        '0' when "0111010011",
        '1' when "0111010100",
        '0' when "0111010101",
        '1' when "0111010110",
        '0' when "0111010111",
        '1' when "0111011000",
        '0' when "0111011001",
        '1' when "0111011010",
        '0' when "0111011011",
        '1' when "0111011100",
        '0' when "0111011101",
        '1' when "0111011110",
        '0' when "0111011111",
        '1' when "0111100000",
        '0' when "0111100001",
        '1' when "0111100010",
        '0' when "0111100011",
        '1' when "0111100100",
        '0' when "0111100101",
        '1' when "0111100110",
        '0' when "0111100111",
        '1' when "0111101000",
        '0' when "0111101001",
        '1' when "0111101010",
        '0' when "0111101011",
        '1' when "0111101100",
        '0' when "0111101101",
        '1' when "0111101110",
        '0' when "0111101111",
        '1' when "0111110000",
        '0' when "0111110001",
        '1' when "0111110010",
        '0' when "0111110011",
        '1' when "0111110100",
        '0' when "0111110101",
        '1' when "0111110110",
        '0' when "0111110111",
        '1' when "0111111000",
        '0' when "0111111001",
        '1' when "0111111010",
        '0' when "0111111011",
        '1' when "0111111100",
        '0' when "0111111101",
        '1' when "0111111110",
        '0' when "0111111111",
        '1' when "1000000000",
        '0' when "1000000001",
        '1' when "1000000010",
        '0' when "1000000011",
        '1' when "1000000100",
        '0' when "1000000101",
        '1' when "1000000110",
        '0' when "1000000111",
        '1' when "1000001000",
        '0' when "1000001001",
        '1' when "1000001010",
        '0' when "1000001011",
        '1' when "1000001100",
        '0' when "1000001101",
        '1' when "1000001110",
        '0' when "1000001111",
        '1' when "1000010000",
        '0' when "1000010001",
        '1' when "1000010010",
        '0' when "1000010011",
        '1' when "1000010100",
        '0' when "1000010101",
        '1' when "1000010110",
        '0' when "1000010111",
        '1' when "1000011000",
        '0' when "1000011001",
        '1' when "1000011010",
        '0' when "1000011011",
        '1' when "1000011100",
        '0' when "1000011101",
        '1' when "1000011110",
        '0' when "1000011111",
        '1' when "1000100000",
        '0' when "1000100001",
        '1' when "1000100010",
        '0' when "1000100011",
        '1' when "1000100100",
        '0' when "1000100101",
        '1' when "1000100110",
        '0' when "1000100111",
        '1' when "1000101000",
        '0' when "1000101001",
        '1' when "1000101010",
        '0' when "1000101011",
        '1' when "1000101100",
        '0' when "1000101101",
        '1' when "1000101110",
        '0' when "1000101111",
        '1' when "1000110000",
        '0' when "1000110001",
        '1' when "1000110010",
        '0' when "1000110011",
        '1' when "1000110100",
        '0' when "1000110101",
        '1' when "1000110110",
        '0' when "1000110111",
        '1' when "1000111000",
        '0' when "1000111001",
        '1' when "1000111010",
        '0' when "1000111011",
        '1' when "1000111100",
        '0' when "1000111101",
        '1' when "1000111110",
        '0' when "1000111111",
        '1' when "1001000000",
        '0' when "1001000001",
        '1' when "1001000010",
        '0' when "1001000011",
        '1' when "1001000100",
        '0' when "1001000101",
        '1' when "1001000110",
        '0' when "1001000111",
        '1' when "1001001000",
        '0' when "1001001001",
        '1' when "1001001010",
        '0' when "1001001011",
        '1' when "1001001100",
        '0' when "1001001101",
        '1' when "1001001110",
        '0' when "1001001111",
        '1' when "1001010000",
        '0' when "1001010001",
        '1' when "1001010010",
        '0' when "1001010011",
        '1' when "1001010100",
        '0' when "1001010101",
        '1' when "1001010110",
        '0' when "1001010111",
        '1' when "1001011000",
        '0' when "1001011001",
        '1' when "1001011010",
        '0' when "1001011011",
        '1' when "1001011100",
        '0' when "1001011101",
        '1' when "1001011110",
        '0' when "1001011111",
        '1' when "1001100000",
        '0' when "1001100001",
        '1' when "1001100010",
        '0' when "1001100011",
        '1' when "1001100100",
        '0' when "1001100101",
        '1' when "1001100110",
        '0' when "1001100111",
        '1' when "1001101000",
        '0' when "1001101001",
        '1' when "1001101010",
        '0' when "1001101011",
        '1' when "1001101100",
        '0' when "1001101101",
        '1' when "1001101110",
        '0' when "1001101111",
        '1' when "1001110000",
        '0' when "1001110001",
        '1' when "1001110010",
        '0' when "1001110011",
        '1' when "1001110100",
        '0' when "1001110101",
        '1' when "1001110110",
        '0' when "1001110111",
        '1' when "1001111000",
        '0' when "1001111001",
        '1' when "1001111010",
        '0' when "1001111011",
        '1' when "1001111100",
        '0' when "1001111101",
        '1' when "1001111110",
        '0' when "1001111111",
        '1' when "1010000000",
        '0' when "1010000001",
        '1' when "1010000010",
        '0' when "1010000011",
        '1' when "1010000100",
        '0' when "1010000101",
        '1' when "1010000110",
        '0' when "1010000111",
        '1' when "1010001000",
        '0' when "1010001001",
        '1' when "1010001010",
        '0' when "1010001011",
        '1' when "1010001100",
        '0' when "1010001101",
        '1' when "1010001110",
        '0' when "1010001111",
        '1' when "1010010000",
        '0' when "1010010001",
        '1' when "1010010010",
        '0' when "1010010011",
        '1' when "1010010100",
        '0' when "1010010101",
        '1' when "1010010110",
        '0' when "1010010111",
        '1' when "1010011000",
        '0' when "1010011001",
        '1' when "1010011010",
        '0' when "1010011011",
        '1' when "1010011100",
        '0' when "1010011101",
        '1' when "1010011110",
        '0' when "1010011111",
        '1' when "1010100000",
        '0' when "1010100001",
        '1' when "1010100010",
        '0' when "1010100011",
        '1' when "1010100100",
        '0' when "1010100101",
        '1' when "1010100110",
        '0' when "1010100111",
        '1' when "1010101000",
        '0' when "1010101001",
        '1' when "1010101010",
        '0' when "1010101011",
        '1' when "1010101100",
        '0' when "1010101101",
        '1' when "1010101110",
        '0' when "1010101111",
        '1' when "1010110000",
        '0' when "1010110001",
        '1' when "1010110010",
        '0' when "1010110011",
        '1' when "1010110100",
        '0' when "1010110101",
        '1' when "1010110110",
        '0' when "1010110111",
        '1' when "1010111000",
        '0' when "1010111001",
        '1' when "1010111010",
        '0' when "1010111011",
        '1' when "1010111100",
        '0' when "1010111101",
        '1' when "1010111110",
        '0' when "1010111111",
        '1' when "1011000000",
        '0' when "1011000001",
        '1' when "1011000010",
        '0' when "1011000011",
        '1' when "1011000100",
        '0' when "1011000101",
        '1' when "1011000110",
        '0' when "1011000111",
        '1' when "1011001000",
        '0' when "1011001001",
        '1' when "1011001010",
        '0' when "1011001011",
        '1' when "1011001100",
        '0' when "1011001101",
        '1' when "1011001110",
        '0' when "1011001111",
        '1' when "1011010000",
        '0' when "1011010001",
        '1' when "1011010010",
        '0' when "1011010011",
        '1' when "1011010100",
        '0' when "1011010101",
        '1' when "1011010110",
        '0' when "1011010111",
        '1' when "1011011000",
        '0' when "1011011001",
        '1' when "1011011010",
        '0' when "1011011011",
        '1' when "1011011100",
        '0' when "1011011101",
        '1' when "1011011110",
        '0' when "1011011111",
        '1' when "1011100000",
        '0' when "1011100001",
        '1' when "1011100010",
        '0' when "1011100011",
        '1' when "1011100100",
        '0' when "1011100101",
        '1' when "1011100110",
        '0' when "1011100111",
        '1' when "1011101000",
        '0' when "1011101001",
        '1' when "1011101010",
        '0' when "1011101011",
        '1' when "1011101100",
        '0' when "1011101101",
        '1' when "1011101110",
        '0' when "1011101111",
        '1' when "1011110000",
        '0' when "1011110001",
        '1' when "1011110010",
        '0' when "1011110011",
        '1' when "1011110100",
        '0' when "1011110101",
        '1' when "1011110110",
        '0' when "1011110111",
        '1' when "1011111000",
        '0' when "1011111001",
        '1' when "1011111010",
        '0' when "1011111011",
        '1' when "1011111100",
        '0' when "1011111101",
        '1' when "1011111110",
        '0' when "1011111111",
        '1' when "1100000000",
        '0' when "1100000001",
        '1' when "1100000010",
        '0' when "1100000011",
        '1' when "1100000100",
        '0' when "1100000101",
        '1' when "1100000110",
        '0' when "1100000111",
        '1' when "1100001000",
        '0' when "1100001001",
        '1' when "1100001010",
        '0' when "1100001011",
        '1' when "1100001100",
        '0' when "1100001101",
        '1' when "1100001110",
        '0' when "1100001111",
        '1' when "1100010000",
        '0' when "1100010001",
        '1' when "1100010010",
        '0' when "1100010011",
        '1' when "1100010100",
        '0' when "1100010101",
        '1' when "1100010110",
        '0' when "1100010111",
        '1' when "1100011000",
        '0' when "1100011001",
        '1' when "1100011010",
        '0' when "1100011011",
        '1' when "1100011100",
        '0' when "1100011101",
        '1' when "1100011110",
        '0' when "1100011111",
        '1' when "1100100000",
        '0' when "1100100001",
        '1' when "1100100010",
        '0' when "1100100011",
        '1' when "1100100100",
        '0' when "1100100101",
        '1' when "1100100110",
        '0' when "1100100111",
        '1' when "1100101000",
        '0' when "1100101001",
        '1' when "1100101010",
        '0' when "1100101011",
        '1' when "1100101100",
        '0' when "1100101101",
        '1' when "1100101110",
        '0' when "1100101111",
        '1' when "1100110000",
        '0' when "1100110001",
        '1' when "1100110010",
        '0' when "1100110011",
        '1' when "1100110100",
        '0' when "1100110101",
        '1' when "1100110110",
        '0' when "1100110111",
        '1' when "1100111000",
        '0' when "1100111001",
        '1' when "1100111010",
        '0' when "1100111011",
        '1' when "1100111100",
        '0' when "1100111101",
        '1' when "1100111110",
        '0' when "1100111111",
        '1' when "1101000000",
        '0' when "1101000001",
        '1' when "1101000010",
        '0' when "1101000011",
        '1' when "1101000100",
        '0' when "1101000101",
        '1' when "1101000110",
        '0' when "1101000111",
        '1' when "1101001000",
        '0' when "1101001001",
        '1' when "1101001010",
        '0' when "1101001011",
        '1' when "1101001100",
        '0' when "1101001101",
        '1' when "1101001110",
        '0' when "1101001111",
        '1' when "1101010000",
        '0' when "1101010001",
        '1' when "1101010010",
        '0' when "1101010011",
        '1' when "1101010100",
        '0' when "1101010101",
        '1' when "1101010110",
        '0' when "1101010111",
        '1' when "1101011000",
        '0' when "1101011001",
        '1' when "1101011010",
        '0' when "1101011011",
        '1' when "1101011100",
        '0' when "1101011101",
        '1' when "1101011110",
        '0' when "1101011111",
        '1' when "1101100000",
        '0' when "1101100001",
        '1' when "1101100010",
        '0' when "1101100011",
        '1' when "1101100100",
        '0' when "1101100101",
        '1' when "1101100110",
        '0' when "1101100111",
        '1' when "1101101000",
        '0' when "1101101001",
        '1' when "1101101010",
        '0' when "1101101011",
        '1' when "1101101100",
        '0' when "1101101101",
        '1' when "1101101110",
        '0' when "1101101111",
        '1' when "1101110000",
        '0' when "1101110001",
        '1' when "1101110010",
        '0' when "1101110011",
        '1' when "1101110100",
        '0' when "1101110101",
        '1' when "1101110110",
        '0' when "1101110111",
        '1' when "1101111000",
        '0' when "1101111001",
        '1' when "1101111010",
        '0' when "1101111011",
        '1' when "1101111100",
        '0' when "1101111101",
        '1' when "1101111110",
        '0' when "1101111111",
        '1' when "1110000000",
        '0' when "1110000001",
        '1' when "1110000010",
        '0' when "1110000011",
        '1' when "1110000100",
        '0' when "1110000101",
        '1' when "1110000110",
        '0' when "1110000111",
        '1' when "1110001000",
        '0' when "1110001001",
        '1' when "1110001010",
        '0' when "1110001011",
        '1' when "1110001100",
        '0' when "1110001101",
        '1' when "1110001110",
        '0' when "1110001111",
        '1' when "1110010000",
        '0' when "1110010001",
        '1' when "1110010010",
        '0' when "1110010011",
        '1' when "1110010100",
        '0' when "1110010101",
        '1' when "1110010110",
        '0' when "1110010111",
        '1' when "1110011000",
        '0' when "1110011001",
        '1' when "1110011010",
        '0' when "1110011011",
        '1' when "1110011100",
        '0' when "1110011101",
        '1' when "1110011110",
        '0' when "1110011111",
        '1' when "1110100000",
        '0' when "1110100001",
        '1' when "1110100010",
        '0' when "1110100011",
        '1' when "1110100100",
        '0' when "1110100101",
        '1' when "1110100110",
        '0' when "1110100111",
        '1' when "1110101000",
        '0' when "1110101001",
        '1' when "1110101010",
        '0' when "1110101011",
        '1' when "1110101100",
        '0' when "1110101101",
        '1' when "1110101110",
        '0' when "1110101111",
        '1' when "1110110000",
        '0' when "1110110001",
        '1' when "1110110010",
        '0' when "1110110011",
        '1' when "1110110100",
        '0' when "1110110101",
        '1' when "1110110110",
        '0' when "1110110111",
        '1' when "1110111000",
        '0' when "1110111001",
        '1' when "1110111010",
        '0' when "1110111011",
        '1' when "1110111100",
        '0' when "1110111101",
        '1' when "1110111110",
        '0' when "1110111111",
        '1' when "1111000000",
        '0' when "1111000001",
        '1' when "1111000010",
        '0' when "1111000011",
        '1' when "1111000100",
        '0' when "1111000101",
        '1' when "1111000110",
        '0' when "1111000111",
        '1' when "1111001000",
        '0' when "1111001001",
        '1' when "1111001010",
        '0' when "1111001011",
        '1' when "1111001100",
        '0' when "1111001101",
        '1' when "1111001110",
        '0' when "1111001111",
        '1' when "1111010000",
        '0' when "1111010001",
        '1' when "1111010010",
        '0' when "1111010011",
        '1' when "1111010100",
        '0' when "1111010101",
        '1' when "1111010110",
        '0' when "1111010111",
        '1' when "1111011000",
        '0' when "1111011001",
        '1' when "1111011010",
        '0' when "1111011011",
        '1' when "1111011100",
        '0' when "1111011101",
        '1' when "1111011110",
        '0' when "1111011111",
        '1' when "1111100000",
        '0' when "1111100001",
        '1' when "1111100010",
        '0' when "1111100011",
        '1' when "1111100100",
        '0' when "1111100101",
        '1' when "1111100110",
        '0' when "1111100111",
        '1' when "1111101000",
        '0' when "1111101001",
        '1' when "1111101010",
        '0' when "1111101011",
        '1' when "1111101100",
        '0' when "1111101101",
        '1' when "1111101110",
        '0' when "1111101111",
        '1' when "1111110000",
        '0' when "1111110001",
        '1' when "1111110010",
        '0' when "1111110011",
        '1' when "1111110100",
        '0' when "1111110101",
        '1' when "1111110110",
        '0' when "1111110111",
        '1' when "1111111000",
        '0' when "1111111001",
        '1' when "1111111010",
        '0' when "1111111011",
        '1' when "1111111100",
        '0' when "1111111101",
        '1' when "1111111110",
        '0' when "1111111111",
        '0' when others;

    -- Truth table for when number is odd
    with concatenatedBits select odd <=
        '0' when "0000000000",
        '1' when "0000000001",
        '0' when "0000000010",
        '1' when "0000000011",
        '0' when "0000000100",
        '1' when "0000000101",
        '0' when "0000000110",
        '1' when "0000000111",
        '0' when "0000001000",
        '1' when "0000001001",
        '0' when "0000001010",
        '1' when "0000001011",
        '0' when "0000001100",
        '1' when "0000001101",
        '0' when "0000001110",
        '1' when "0000001111",
        '0' when "0000010000",
        '1' when "0000010001",
        '0' when "0000010010",
        '1' when "0000010011",
        '0' when "0000010100",
        '1' when "0000010101",
        '0' when "0000010110",
        '1' when "0000010111",
        '0' when "0000011000",
        '1' when "0000011001",
        '0' when "0000011010",
        '1' when "0000011011",
        '0' when "0000011100",
        '1' when "0000011101",
        '0' when "0000011110",
        '1' when "0000011111",
        '0' when "0000100000",
        '1' when "0000100001",
        '0' when "0000100010",
        '1' when "0000100011",
        '0' when "0000100100",
        '1' when "0000100101",
        '0' when "0000100110",
        '1' when "0000100111",
        '0' when "0000101000",
        '1' when "0000101001",
        '0' when "0000101010",
        '1' when "0000101011",
        '0' when "0000101100",
        '1' when "0000101101",
        '0' when "0000101110",
        '1' when "0000101111",
        '0' when "0000110000",
        '1' when "0000110001",
        '0' when "0000110010",
        '1' when "0000110011",
        '0' when "0000110100",
        '1' when "0000110101",
        '0' when "0000110110",
        '1' when "0000110111",
        '0' when "0000111000",
        '1' when "0000111001",
        '0' when "0000111010",
        '1' when "0000111011",
        '0' when "0000111100",
        '1' when "0000111101",
        '0' when "0000111110",
        '1' when "0000111111",
        '0' when "0001000000",
        '1' when "0001000001",
        '0' when "0001000010",
        '1' when "0001000011",
        '0' when "0001000100",
        '1' when "0001000101",
        '0' when "0001000110",
        '1' when "0001000111",
        '0' when "0001001000",
        '1' when "0001001001",
        '0' when "0001001010",
        '1' when "0001001011",
        '0' when "0001001100",
        '1' when "0001001101",
        '0' when "0001001110",
        '1' when "0001001111",
        '0' when "0001010000",
        '1' when "0001010001",
        '0' when "0001010010",
        '1' when "0001010011",
        '0' when "0001010100",
        '1' when "0001010101",
        '0' when "0001010110",
        '1' when "0001010111",
        '0' when "0001011000",
        '1' when "0001011001",
        '0' when "0001011010",
        '1' when "0001011011",
        '0' when "0001011100",
        '1' when "0001011101",
        '0' when "0001011110",
        '1' when "0001011111",
        '0' when "0001100000",
        '1' when "0001100001",
        '0' when "0001100010",
        '1' when "0001100011",
        '0' when "0001100100",
        '1' when "0001100101",
        '0' when "0001100110",
        '1' when "0001100111",
        '0' when "0001101000",
        '1' when "0001101001",
        '0' when "0001101010",
        '1' when "0001101011",
        '0' when "0001101100",
        '1' when "0001101101",
        '0' when "0001101110",
        '1' when "0001101111",
        '0' when "0001110000",
        '1' when "0001110001",
        '0' when "0001110010",
        '1' when "0001110011",
        '0' when "0001110100",
        '1' when "0001110101",
        '0' when "0001110110",
        '1' when "0001110111",
        '0' when "0001111000",
        '1' when "0001111001",
        '0' when "0001111010",
        '1' when "0001111011",
        '0' when "0001111100",
        '1' when "0001111101",
        '0' when "0001111110",
        '1' when "0001111111",
        '0' when "0010000000",
        '1' when "0010000001",
        '0' when "0010000010",
        '1' when "0010000011",
        '0' when "0010000100",
        '1' when "0010000101",
        '0' when "0010000110",
        '1' when "0010000111",
        '0' when "0010001000",
        '1' when "0010001001",
        '0' when "0010001010",
        '1' when "0010001011",
        '0' when "0010001100",
        '1' when "0010001101",
        '0' when "0010001110",
        '1' when "0010001111",
        '0' when "0010010000",
        '1' when "0010010001",
        '0' when "0010010010",
        '1' when "0010010011",
        '0' when "0010010100",
        '1' when "0010010101",
        '0' when "0010010110",
        '1' when "0010010111",
        '0' when "0010011000",
        '1' when "0010011001",
        '0' when "0010011010",
        '1' when "0010011011",
        '0' when "0010011100",
        '1' when "0010011101",
        '0' when "0010011110",
        '1' when "0010011111",
        '0' when "0010100000",
        '1' when "0010100001",
        '0' when "0010100010",
        '1' when "0010100011",
        '0' when "0010100100",
        '1' when "0010100101",
        '0' when "0010100110",
        '1' when "0010100111",
        '0' when "0010101000",
        '1' when "0010101001",
        '0' when "0010101010",
        '1' when "0010101011",
        '0' when "0010101100",
        '1' when "0010101101",
        '0' when "0010101110",
        '1' when "0010101111",
        '0' when "0010110000",
        '1' when "0010110001",
        '0' when "0010110010",
        '1' when "0010110011",
        '0' when "0010110100",
        '1' when "0010110101",
        '0' when "0010110110",
        '1' when "0010110111",
        '0' when "0010111000",
        '1' when "0010111001",
        '0' when "0010111010",
        '1' when "0010111011",
        '0' when "0010111100",
        '1' when "0010111101",
        '0' when "0010111110",
        '1' when "0010111111",
        '0' when "0011000000",
        '1' when "0011000001",
        '0' when "0011000010",
        '1' when "0011000011",
        '0' when "0011000100",
        '1' when "0011000101",
        '0' when "0011000110",
        '1' when "0011000111",
        '0' when "0011001000",
        '1' when "0011001001",
        '0' when "0011001010",
        '1' when "0011001011",
        '0' when "0011001100",
        '1' when "0011001101",
        '0' when "0011001110",
        '1' when "0011001111",
        '0' when "0011010000",
        '1' when "0011010001",
        '0' when "0011010010",
        '1' when "0011010011",
        '0' when "0011010100",
        '1' when "0011010101",
        '0' when "0011010110",
        '1' when "0011010111",
        '0' when "0011011000",
        '1' when "0011011001",
        '0' when "0011011010",
        '1' when "0011011011",
        '0' when "0011011100",
        '1' when "0011011101",
        '0' when "0011011110",
        '1' when "0011011111",
        '0' when "0011100000",
        '1' when "0011100001",
        '0' when "0011100010",
        '1' when "0011100011",
        '0' when "0011100100",
        '1' when "0011100101",
        '0' when "0011100110",
        '1' when "0011100111",
        '0' when "0011101000",
        '1' when "0011101001",
        '0' when "0011101010",
        '1' when "0011101011",
        '0' when "0011101100",
        '1' when "0011101101",
        '0' when "0011101110",
        '1' when "0011101111",
        '0' when "0011110000",
        '1' when "0011110001",
        '0' when "0011110010",
        '1' when "0011110011",
        '0' when "0011110100",
        '1' when "0011110101",
        '0' when "0011110110",
        '1' when "0011110111",
        '0' when "0011111000",
        '1' when "0011111001",
        '0' when "0011111010",
        '1' when "0011111011",
        '0' when "0011111100",
        '1' when "0011111101",
        '0' when "0011111110",
        '1' when "0011111111",
        '0' when "0100000000",
        '1' when "0100000001",
        '0' when "0100000010",
        '1' when "0100000011",
        '0' when "0100000100",
        '1' when "0100000101",
        '0' when "0100000110",
        '1' when "0100000111",
        '0' when "0100001000",
        '1' when "0100001001",
        '0' when "0100001010",
        '1' when "0100001011",
        '0' when "0100001100",
        '1' when "0100001101",
        '0' when "0100001110",
        '1' when "0100001111",
        '0' when "0100010000",
        '1' when "0100010001",
        '0' when "0100010010",
        '1' when "0100010011",
        '0' when "0100010100",
        '1' when "0100010101",
        '0' when "0100010110",
        '1' when "0100010111",
        '0' when "0100011000",
        '1' when "0100011001",
        '0' when "0100011010",
        '1' when "0100011011",
        '0' when "0100011100",
        '1' when "0100011101",
        '0' when "0100011110",
        '1' when "0100011111",
        '0' when "0100100000",
        '1' when "0100100001",
        '0' when "0100100010",
        '1' when "0100100011",
        '0' when "0100100100",
        '1' when "0100100101",
        '0' when "0100100110",
        '1' when "0100100111",
        '0' when "0100101000",
        '1' when "0100101001",
        '0' when "0100101010",
        '1' when "0100101011",
        '0' when "0100101100",
        '1' when "0100101101",
        '0' when "0100101110",
        '1' when "0100101111",
        '0' when "0100110000",
        '1' when "0100110001",
        '0' when "0100110010",
        '1' when "0100110011",
        '0' when "0100110100",
        '1' when "0100110101",
        '0' when "0100110110",
        '1' when "0100110111",
        '0' when "0100111000",
        '1' when "0100111001",
        '0' when "0100111010",
        '1' when "0100111011",
        '0' when "0100111100",
        '1' when "0100111101",
        '0' when "0100111110",
        '1' when "0100111111",
        '0' when "0101000000",
        '1' when "0101000001",
        '0' when "0101000010",
        '1' when "0101000011",
        '0' when "0101000100",
        '1' when "0101000101",
        '0' when "0101000110",
        '1' when "0101000111",
        '0' when "0101001000",
        '1' when "0101001001",
        '0' when "0101001010",
        '1' when "0101001011",
        '0' when "0101001100",
        '1' when "0101001101",
        '0' when "0101001110",
        '1' when "0101001111",
        '0' when "0101010000",
        '1' when "0101010001",
        '0' when "0101010010",
        '1' when "0101010011",
        '0' when "0101010100",
        '1' when "0101010101",
        '0' when "0101010110",
        '1' when "0101010111",
        '0' when "0101011000",
        '1' when "0101011001",
        '0' when "0101011010",
        '1' when "0101011011",
        '0' when "0101011100",
        '1' when "0101011101",
        '0' when "0101011110",
        '1' when "0101011111",
        '0' when "0101100000",
        '1' when "0101100001",
        '0' when "0101100010",
        '1' when "0101100011",
        '0' when "0101100100",
        '1' when "0101100101",
        '0' when "0101100110",
        '1' when "0101100111",
        '0' when "0101101000",
        '1' when "0101101001",
        '0' when "0101101010",
        '1' when "0101101011",
        '0' when "0101101100",
        '1' when "0101101101",
        '0' when "0101101110",
        '1' when "0101101111",
        '0' when "0101110000",
        '1' when "0101110001",
        '0' when "0101110010",
        '1' when "0101110011",
        '0' when "0101110100",
        '1' when "0101110101",
        '0' when "0101110110",
        '1' when "0101110111",
        '0' when "0101111000",
        '1' when "0101111001",
        '0' when "0101111010",
        '1' when "0101111011",
        '0' when "0101111100",
        '1' when "0101111101",
        '0' when "0101111110",
        '1' when "0101111111",
        '0' when "0110000000",
        '1' when "0110000001",
        '0' when "0110000010",
        '1' when "0110000011",
        '0' when "0110000100",
        '1' when "0110000101",
        '0' when "0110000110",
        '1' when "0110000111",
        '0' when "0110001000",
        '1' when "0110001001",
        '0' when "0110001010",
        '1' when "0110001011",
        '0' when "0110001100",
        '1' when "0110001101",
        '0' when "0110001110",
        '1' when "0110001111",
        '0' when "0110010000",
        '1' when "0110010001",
        '0' when "0110010010",
        '1' when "0110010011",
        '0' when "0110010100",
        '1' when "0110010101",
        '0' when "0110010110",
        '1' when "0110010111",
        '0' when "0110011000",
        '1' when "0110011001",
        '0' when "0110011010",
        '1' when "0110011011",
        '0' when "0110011100",
        '1' when "0110011101",
        '0' when "0110011110",
        '1' when "0110011111",
        '0' when "0110100000",
        '1' when "0110100001",
        '0' when "0110100010",
        '1' when "0110100011",
        '0' when "0110100100",
        '1' when "0110100101",
        '0' when "0110100110",
        '1' when "0110100111",
        '0' when "0110101000",
        '1' when "0110101001",
        '0' when "0110101010",
        '1' when "0110101011",
        '0' when "0110101100",
        '1' when "0110101101",
        '0' when "0110101110",
        '1' when "0110101111",
        '0' when "0110110000",
        '1' when "0110110001",
        '0' when "0110110010",
        '1' when "0110110011",
        '0' when "0110110100",
        '1' when "0110110101",
        '0' when "0110110110",
        '1' when "0110110111",
        '0' when "0110111000",
        '1' when "0110111001",
        '0' when "0110111010",
        '1' when "0110111011",
        '0' when "0110111100",
        '1' when "0110111101",
        '0' when "0110111110",
        '1' when "0110111111",
        '0' when "0111000000",
        '1' when "0111000001",
        '0' when "0111000010",
        '1' when "0111000011",
        '0' when "0111000100",
        '1' when "0111000101",
        '0' when "0111000110",
        '1' when "0111000111",
        '0' when "0111001000",
        '1' when "0111001001",
        '0' when "0111001010",
        '1' when "0111001011",
        '0' when "0111001100",
        '1' when "0111001101",
        '0' when "0111001110",
        '1' when "0111001111",
        '0' when "0111010000",
        '1' when "0111010001",
        '0' when "0111010010",
        '1' when "0111010011",
        '0' when "0111010100",
        '1' when "0111010101",
        '0' when "0111010110",
        '1' when "0111010111",
        '0' when "0111011000",
        '1' when "0111011001",
        '0' when "0111011010",
        '1' when "0111011011",
        '0' when "0111011100",
        '1' when "0111011101",
        '0' when "0111011110",
        '1' when "0111011111",
        '0' when "0111100000",
        '1' when "0111100001",
        '0' when "0111100010",
        '1' when "0111100011",
        '0' when "0111100100",
        '1' when "0111100101",
        '0' when "0111100110",
        '1' when "0111100111",
        '0' when "0111101000",
        '1' when "0111101001",
        '0' when "0111101010",
        '1' when "0111101011",
        '0' when "0111101100",
        '1' when "0111101101",
        '0' when "0111101110",
        '1' when "0111101111",
        '0' when "0111110000",
        '1' when "0111110001",
        '0' when "0111110010",
        '1' when "0111110011",
        '0' when "0111110100",
        '1' when "0111110101",
        '0' when "0111110110",
        '1' when "0111110111",
        '0' when "0111111000",
        '1' when "0111111001",
        '0' when "0111111010",
        '1' when "0111111011",
        '0' when "0111111100",
        '1' when "0111111101",
        '0' when "0111111110",
        '1' when "0111111111",
        '0' when "1000000000",
        '1' when "1000000001",
        '0' when "1000000010",
        '1' when "1000000011",
        '0' when "1000000100",
        '1' when "1000000101",
        '0' when "1000000110",
        '1' when "1000000111",
        '0' when "1000001000",
        '1' when "1000001001",
        '0' when "1000001010",
        '1' when "1000001011",
        '0' when "1000001100",
        '1' when "1000001101",
        '0' when "1000001110",
        '1' when "1000001111",
        '0' when "1000010000",
        '1' when "1000010001",
        '0' when "1000010010",
        '1' when "1000010011",
        '0' when "1000010100",
        '1' when "1000010101",
        '0' when "1000010110",
        '1' when "1000010111",
        '0' when "1000011000",
        '1' when "1000011001",
        '0' when "1000011010",
        '1' when "1000011011",
        '0' when "1000011100",
        '1' when "1000011101",
        '0' when "1000011110",
        '1' when "1000011111",
        '0' when "1000100000",
        '1' when "1000100001",
        '0' when "1000100010",
        '1' when "1000100011",
        '0' when "1000100100",
        '1' when "1000100101",
        '0' when "1000100110",
        '1' when "1000100111",
        '0' when "1000101000",
        '1' when "1000101001",
        '0' when "1000101010",
        '1' when "1000101011",
        '0' when "1000101100",
        '1' when "1000101101",
        '0' when "1000101110",
        '1' when "1000101111",
        '0' when "1000110000",
        '1' when "1000110001",
        '0' when "1000110010",
        '1' when "1000110011",
        '0' when "1000110100",
        '1' when "1000110101",
        '0' when "1000110110",
        '1' when "1000110111",
        '0' when "1000111000",
        '1' when "1000111001",
        '0' when "1000111010",
        '1' when "1000111011",
        '0' when "1000111100",
        '1' when "1000111101",
        '0' when "1000111110",
        '1' when "1000111111",
        '0' when "1001000000",
        '1' when "1001000001",
        '0' when "1001000010",
        '1' when "1001000011",
        '0' when "1001000100",
        '1' when "1001000101",
        '0' when "1001000110",
        '1' when "1001000111",
        '0' when "1001001000",
        '1' when "1001001001",
        '0' when "1001001010",
        '1' when "1001001011",
        '0' when "1001001100",
        '1' when "1001001101",
        '0' when "1001001110",
        '1' when "1001001111",
        '0' when "1001010000",
        '1' when "1001010001",
        '0' when "1001010010",
        '1' when "1001010011",
        '0' when "1001010100",
        '1' when "1001010101",
        '0' when "1001010110",
        '1' when "1001010111",
        '0' when "1001011000",
        '1' when "1001011001",
        '0' when "1001011010",
        '1' when "1001011011",
        '0' when "1001011100",
        '1' when "1001011101",
        '0' when "1001011110",
        '1' when "1001011111",
        '0' when "1001100000",
        '1' when "1001100001",
        '0' when "1001100010",
        '1' when "1001100011",
        '0' when "1001100100",
        '1' when "1001100101",
        '0' when "1001100110",
        '1' when "1001100111",
        '0' when "1001101000",
        '1' when "1001101001",
        '0' when "1001101010",
        '1' when "1001101011",
        '0' when "1001101100",
        '1' when "1001101101",
        '0' when "1001101110",
        '1' when "1001101111",
        '0' when "1001110000",
        '1' when "1001110001",
        '0' when "1001110010",
        '1' when "1001110011",
        '0' when "1001110100",
        '1' when "1001110101",
        '0' when "1001110110",
        '1' when "1001110111",
        '0' when "1001111000",
        '1' when "1001111001",
        '0' when "1001111010",
        '1' when "1001111011",
        '0' when "1001111100",
        '1' when "1001111101",
        '0' when "1001111110",
        '1' when "1001111111",
        '0' when "1010000000",
        '1' when "1010000001",
        '0' when "1010000010",
        '1' when "1010000011",
        '0' when "1010000100",
        '1' when "1010000101",
        '0' when "1010000110",
        '1' when "1010000111",
        '0' when "1010001000",
        '1' when "1010001001",
        '0' when "1010001010",
        '1' when "1010001011",
        '0' when "1010001100",
        '1' when "1010001101",
        '0' when "1010001110",
        '1' when "1010001111",
        '0' when "1010010000",
        '1' when "1010010001",
        '0' when "1010010010",
        '1' when "1010010011",
        '0' when "1010010100",
        '1' when "1010010101",
        '0' when "1010010110",
        '1' when "1010010111",
        '0' when "1010011000",
        '1' when "1010011001",
        '0' when "1010011010",
        '1' when "1010011011",
        '0' when "1010011100",
        '1' when "1010011101",
        '0' when "1010011110",
        '1' when "1010011111",
        '0' when "1010100000",
        '1' when "1010100001",
        '0' when "1010100010",
        '1' when "1010100011",
        '0' when "1010100100",
        '1' when "1010100101",
        '0' when "1010100110",
        '1' when "1010100111",
        '0' when "1010101000",
        '1' when "1010101001",
        '0' when "1010101010",
        '1' when "1010101011",
        '0' when "1010101100",
        '1' when "1010101101",
        '0' when "1010101110",
        '1' when "1010101111",
        '0' when "1010110000",
        '1' when "1010110001",
        '0' when "1010110010",
        '1' when "1010110011",
        '0' when "1010110100",
        '1' when "1010110101",
        '0' when "1010110110",
        '1' when "1010110111",
        '0' when "1010111000",
        '1' when "1010111001",
        '0' when "1010111010",
        '1' when "1010111011",
        '0' when "1010111100",
        '1' when "1010111101",
        '0' when "1010111110",
        '1' when "1010111111",
        '0' when "1011000000",
        '1' when "1011000001",
        '0' when "1011000010",
        '1' when "1011000011",
        '0' when "1011000100",
        '1' when "1011000101",
        '0' when "1011000110",
        '1' when "1011000111",
        '0' when "1011001000",
        '1' when "1011001001",
        '0' when "1011001010",
        '1' when "1011001011",
        '0' when "1011001100",
        '1' when "1011001101",
        '0' when "1011001110",
        '1' when "1011001111",
        '0' when "1011010000",
        '1' when "1011010001",
        '0' when "1011010010",
        '1' when "1011010011",
        '0' when "1011010100",
        '1' when "1011010101",
        '0' when "1011010110",
        '1' when "1011010111",
        '0' when "1011011000",
        '1' when "1011011001",
        '0' when "1011011010",
        '1' when "1011011011",
        '0' when "1011011100",
        '1' when "1011011101",
        '0' when "1011011110",
        '1' when "1011011111",
        '0' when "1011100000",
        '1' when "1011100001",
        '0' when "1011100010",
        '1' when "1011100011",
        '0' when "1011100100",
        '1' when "1011100101",
        '0' when "1011100110",
        '1' when "1011100111",
        '0' when "1011101000",
        '1' when "1011101001",
        '0' when "1011101010",
        '1' when "1011101011",
        '0' when "1011101100",
        '1' when "1011101101",
        '0' when "1011101110",
        '1' when "1011101111",
        '0' when "1011110000",
        '1' when "1011110001",
        '0' when "1011110010",
        '1' when "1011110011",
        '0' when "1011110100",
        '1' when "1011110101",
        '0' when "1011110110",
        '1' when "1011110111",
        '0' when "1011111000",
        '1' when "1011111001",
        '0' when "1011111010",
        '1' when "1011111011",
        '0' when "1011111100",
        '1' when "1011111101",
        '0' when "1011111110",
        '1' when "1011111111",
        '0' when "1100000000",
        '1' when "1100000001",
        '0' when "1100000010",
        '1' when "1100000011",
        '0' when "1100000100",
        '1' when "1100000101",
        '0' when "1100000110",
        '1' when "1100000111",
        '0' when "1100001000",
        '1' when "1100001001",
        '0' when "1100001010",
        '1' when "1100001011",
        '0' when "1100001100",
        '1' when "1100001101",
        '0' when "1100001110",
        '1' when "1100001111",
        '0' when "1100010000",
        '1' when "1100010001",
        '0' when "1100010010",
        '1' when "1100010011",
        '0' when "1100010100",
        '1' when "1100010101",
        '0' when "1100010110",
        '1' when "1100010111",
        '0' when "1100011000",
        '1' when "1100011001",
        '0' when "1100011010",
        '1' when "1100011011",
        '0' when "1100011100",
        '1' when "1100011101",
        '0' when "1100011110",
        '1' when "1100011111",
        '0' when "1100100000",
        '1' when "1100100001",
        '0' when "1100100010",
        '1' when "1100100011",
        '0' when "1100100100",
        '1' when "1100100101",
        '0' when "1100100110",
        '1' when "1100100111",
        '0' when "1100101000",
        '1' when "1100101001",
        '0' when "1100101010",
        '1' when "1100101011",
        '0' when "1100101100",
        '1' when "1100101101",
        '0' when "1100101110",
        '1' when "1100101111",
        '0' when "1100110000",
        '1' when "1100110001",
        '0' when "1100110010",
        '1' when "1100110011",
        '0' when "1100110100",
        '1' when "1100110101",
        '0' when "1100110110",
        '1' when "1100110111",
        '0' when "1100111000",
        '1' when "1100111001",
        '0' when "1100111010",
        '1' when "1100111011",
        '0' when "1100111100",
        '1' when "1100111101",
        '0' when "1100111110",
        '1' when "1100111111",
        '0' when "1101000000",
        '1' when "1101000001",
        '0' when "1101000010",
        '1' when "1101000011",
        '0' when "1101000100",
        '1' when "1101000101",
        '0' when "1101000110",
        '1' when "1101000111",
        '0' when "1101001000",
        '1' when "1101001001",
        '0' when "1101001010",
        '1' when "1101001011",
        '0' when "1101001100",
        '1' when "1101001101",
        '0' when "1101001110",
        '1' when "1101001111",
        '0' when "1101010000",
        '1' when "1101010001",
        '0' when "1101010010",
        '1' when "1101010011",
        '0' when "1101010100",
        '1' when "1101010101",
        '0' when "1101010110",
        '1' when "1101010111",
        '0' when "1101011000",
        '1' when "1101011001",
        '0' when "1101011010",
        '1' when "1101011011",
        '0' when "1101011100",
        '1' when "1101011101",
        '0' when "1101011110",
        '1' when "1101011111",
        '0' when "1101100000",
        '1' when "1101100001",
        '0' when "1101100010",
        '1' when "1101100011",
        '0' when "1101100100",
        '1' when "1101100101",
        '0' when "1101100110",
        '1' when "1101100111",
        '0' when "1101101000",
        '1' when "1101101001",
        '0' when "1101101010",
        '1' when "1101101011",
        '0' when "1101101100",
        '1' when "1101101101",
        '0' when "1101101110",
        '1' when "1101101111",
        '0' when "1101110000",
        '1' when "1101110001",
        '0' when "1101110010",
        '1' when "1101110011",
        '0' when "1101110100",
        '1' when "1101110101",
        '0' when "1101110110",
        '1' when "1101110111",
        '0' when "1101111000",
        '1' when "1101111001",
        '0' when "1101111010",
        '1' when "1101111011",
        '0' when "1101111100",
        '1' when "1101111101",
        '0' when "1101111110",
        '1' when "1101111111",
        '0' when "1110000000",
        '1' when "1110000001",
        '0' when "1110000010",
        '1' when "1110000011",
        '0' when "1110000100",
        '1' when "1110000101",
        '0' when "1110000110",
        '1' when "1110000111",
        '0' when "1110001000",
        '1' when "1110001001",
        '0' when "1110001010",
        '1' when "1110001011",
        '0' when "1110001100",
        '1' when "1110001101",
        '0' when "1110001110",
        '1' when "1110001111",
        '0' when "1110010000",
        '1' when "1110010001",
        '0' when "1110010010",
        '1' when "1110010011",
        '0' when "1110010100",
        '1' when "1110010101",
        '0' when "1110010110",
        '1' when "1110010111",
        '0' when "1110011000",
        '1' when "1110011001",
        '0' when "1110011010",
        '1' when "1110011011",
        '0' when "1110011100",
        '1' when "1110011101",
        '0' when "1110011110",
        '1' when "1110011111",
        '0' when "1110100000",
        '1' when "1110100001",
        '0' when "1110100010",
        '1' when "1110100011",
        '0' when "1110100100",
        '1' when "1110100101",
        '0' when "1110100110",
        '1' when "1110100111",
        '0' when "1110101000",
        '1' when "1110101001",
        '0' when "1110101010",
        '1' when "1110101011",
        '0' when "1110101100",
        '1' when "1110101101",
        '0' when "1110101110",
        '1' when "1110101111",
        '0' when "1110110000",
        '1' when "1110110001",
        '0' when "1110110010",
        '1' when "1110110011",
        '0' when "1110110100",
        '1' when "1110110101",
        '0' when "1110110110",
        '1' when "1110110111",
        '0' when "1110111000",
        '1' when "1110111001",
        '0' when "1110111010",
        '1' when "1110111011",
        '0' when "1110111100",
        '1' when "1110111101",
        '0' when "1110111110",
        '1' when "1110111111",
        '0' when "1111000000",
        '1' when "1111000001",
        '0' when "1111000010",
        '1' when "1111000011",
        '0' when "1111000100",
        '1' when "1111000101",
        '0' when "1111000110",
        '1' when "1111000111",
        '0' when "1111001000",
        '1' when "1111001001",
        '0' when "1111001010",
        '1' when "1111001011",
        '0' when "1111001100",
        '1' when "1111001101",
        '0' when "1111001110",
        '1' when "1111001111",
        '0' when "1111010000",
        '1' when "1111010001",
        '0' when "1111010010",
        '1' when "1111010011",
        '0' when "1111010100",
        '1' when "1111010101",
        '0' when "1111010110",
        '1' when "1111010111",
        '0' when "1111011000",
        '1' when "1111011001",
        '0' when "1111011010",
        '1' when "1111011011",
        '0' when "1111011100",
        '1' when "1111011101",
        '0' when "1111011110",
        '1' when "1111011111",
        '0' when "1111100000",
        '1' when "1111100001",
        '0' when "1111100010",
        '1' when "1111100011",
        '0' when "1111100100",
        '1' when "1111100101",
        '0' when "1111100110",
        '1' when "1111100111",
        '0' when "1111101000",
        '1' when "1111101001",
        '0' when "1111101010",
        '1' when "1111101011",
        '0' when "1111101100",
        '1' when "1111101101",
        '0' when "1111101110",
        '1' when "1111101111",
        '0' when "1111110000",
        '1' when "1111110001",
        '0' when "1111110010",
        '1' when "1111110011",
        '0' when "1111110100",
        '1' when "1111110101",
        '0' when "1111110110",
        '1' when "1111110111",
        '0' when "1111111000",
        '1' when "1111111001",
        '0' when "1111111010",
        '1' when "1111111011",
        '0' when "1111111100",
        '1' when "1111111101",
        '0' when "1111111110",
        '1' when "1111111111",
        '0' when others;
end tellMeEvenOdd;

-- Thanks for using my library, hope you have memory for it!!
-- (The speeds are theoretically massive, memory is not an issue)